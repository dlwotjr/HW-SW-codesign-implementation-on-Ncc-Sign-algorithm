`timescale 1ns/10ps
`define A #0
